class ahb_seq_clock_glitch extends uvm_sequence #(ahb_seq_item);
  function new(string name = "ahb_seq_clock_glitch");
    super.new(name);
  endfunction

  virtual task body();
    ahb_seq_item item = ahb_seq_item::type_id::create("glitch_item");
    item.addr   = 32'h3A0;
    item.write  = 1;
    item.size   = 3'b010;
    item.burst  = 3'b000;
    item.length = 4;
    item.wdata  = 32'hF00DBABE;
    start_item(item);
    finish_item(item);
    // TB clock overrides during transaction
  endtask

  `uvm_object_utils(ahb_seq_clock_glitch)
endclass

class ahb_test_clock_glitch extends ahb_base_test;
  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  virtual task run_phase(uvm_phase phase);
    phase.raise_objection(this);
    ahb_seq_clock_glitch seq = ahb_seq_clock_glitch::type_id::create("glitch_seq");
    seq.start(env.agent.seqr);
    // Add clock pulse or skip using TB clock thread
    #200ns;
    phase.drop_objection(this);
  endtask

  `uvm_component_utils(ahb_test_clock_glitch)
endclass